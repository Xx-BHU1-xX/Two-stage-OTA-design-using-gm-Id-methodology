.lib "/home/bhuvan/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt
xm1  net-_m1-pad1_ net-_m1-pad2_ gnd gnd sky130_fd_pr__pfet_01v8 W=1 L=0.15
v2 gnd net-_m1-pad1_  dc 1.7
v1 gnd net-_m1-pad2_  dc 1.2
.op
.control
let idval = unitvec(171)
let gmval = unitvec(171)
let gdsval = unitvec(171)
let start = 0
let stop = 1.71
let delta = 0.01
let c = start
while c le stop
alter v1 c
run
let idval[c*100] = @m.xm1.msky130_fd_pr__pfet_01v8[id]
let gmval[c*100] = @m.xm1.msky130_fd_pr__pfet_01v8[gm]
let gdsval[c*100] = @m.xm1.msky130_fd_pr__pfet_01v8[gds]
let c = c + delta
end
setplot new
compose xx start=0 stop=1.7 step=0.01
let idp = idval
let gdsp = gdsval
let gmp = gmval
display
.endc
.end
